
module gem_pad_to_csc_hs_lut(

   input          clock,
   input          wen, // write enable
   input  [7:0]   w_adr, // write address
   input  [7:0]   w_data, // write data

   input          renodd,
   input          reneven,

   input  [7:0]   me1a_r_adr1, 
   output [7:0]   me1a_r_data1, 
   input  [7:0]   me1a_r_adr2, 
   output [7:0]   me1a_r_data2, 
   input  [7:0]   me1b_r_adr1, 
   output [7:0]   me1b_r_data1, 
   input  [7:0]   me1b_r_adr2, 
   output [7:0]   me1b_r_data2 


);


reg [7:0] me1a_r_data1_reg, me1a_r_data2_reg, me1b_r_data1_reg, me1b_r_data2_reg;

always @(posedge clock) begin
    if (wen)   begin
        gem_pad_to_csc_hs_me1a_odd [w_adr] <= w_data; //dump write rom
        gem_pad_to_csc_hs_me1a_even[w_adr] <= w_data;
        gem_pad_to_csc_hs_me1b_odd [w_adr] <= w_data;
        gem_pad_to_csc_hs_me1b_even[w_adr] <= w_data;
    end

    if (renodd)   begin
        me1a_r_data1_reg <= gem_pad_to_csc_hs_me1a_odd[me1a_r_adr1];
        me1a_r_data2_reg <= gem_pad_to_csc_hs_me1a_odd[me1a_r_adr2];
        me1b_r_data1_reg <= gem_pad_to_csc_hs_me1b_odd[me1b_r_adr1];
        me1b_r_data2_reg <= gem_pad_to_csc_hs_me1b_odd[me1b_r_adr2];
    end
    else if (reneven)  begin
        me1a_r_data1_reg <= gem_pad_to_csc_hs_me1a_even[me1a_r_adr1];
        me1a_r_data2_reg <= gem_pad_to_csc_hs_me1a_even[me1a_r_adr2];
        me1b_r_data1_reg <= gem_pad_to_csc_hs_me1b_even[me1b_r_adr1];
        me1b_r_data2_reg <= gem_pad_to_csc_hs_me1b_even[me1b_r_adr2];
    end
end

assign me1a_r_data1 = me1a_r_data1_reg;
assign me1a_r_data2 = me1a_r_data2_reg;
assign me1b_r_data1 = me1b_r_data1_reg;
assign me1b_r_data2 = me1b_r_data2_reg;


reg [ 7:0] gem_pad_to_csc_hs_me1b_odd [191:0];
reg [ 7:0] gem_pad_to_csc_hs_me1b_even [191:0];
reg [ 7:0] gem_pad_to_csc_hs_me1a_odd [191:0];
reg [ 7:0] gem_pad_to_csc_hs_me1a_even [191:0];



  initial begin
	gem_pad_to_csc_hs_me1b_odd[  0]     =   8'd123;
	gem_pad_to_csc_hs_me1b_odd[  1]     =   8'd123;
	gem_pad_to_csc_hs_me1b_odd[  2]     =   8'd122;
	gem_pad_to_csc_hs_me1b_odd[  3]     =   8'd121;
	gem_pad_to_csc_hs_me1b_odd[  4]     =   8'd121;
	gem_pad_to_csc_hs_me1b_odd[  5]     =   8'd120;
	gem_pad_to_csc_hs_me1b_odd[  6]     =   8'd119;
	gem_pad_to_csc_hs_me1b_odd[  7]     =   8'd119;
	gem_pad_to_csc_hs_me1b_odd[  8]     =   8'd118;
	gem_pad_to_csc_hs_me1b_odd[  9]     =   8'd118;
	gem_pad_to_csc_hs_me1b_odd[ 10]     =   8'd117;
	gem_pad_to_csc_hs_me1b_odd[ 11]     =   8'd116;
	gem_pad_to_csc_hs_me1b_odd[ 12]     =   8'd116;
	gem_pad_to_csc_hs_me1b_odd[ 13]     =   8'd115;
	gem_pad_to_csc_hs_me1b_odd[ 14]     =   8'd114;
	gem_pad_to_csc_hs_me1b_odd[ 15]     =   8'd114;
	gem_pad_to_csc_hs_me1b_odd[ 16]     =   8'd113;
	gem_pad_to_csc_hs_me1b_odd[ 17]     =   8'd113;
	gem_pad_to_csc_hs_me1b_odd[ 18]     =   8'd112;
	gem_pad_to_csc_hs_me1b_odd[ 19]     =   8'd111;
	gem_pad_to_csc_hs_me1b_odd[ 20]     =   8'd111;
	gem_pad_to_csc_hs_me1b_odd[ 21]     =   8'd110;
	gem_pad_to_csc_hs_me1b_odd[ 22]     =   8'd110;
	gem_pad_to_csc_hs_me1b_odd[ 23]     =   8'd109;
	gem_pad_to_csc_hs_me1b_odd[ 24]     =   8'd108;
	gem_pad_to_csc_hs_me1b_odd[ 25]     =   8'd108;
	gem_pad_to_csc_hs_me1b_odd[ 26]     =   8'd107;
	gem_pad_to_csc_hs_me1b_odd[ 27]     =   8'd106;
	gem_pad_to_csc_hs_me1b_odd[ 28]     =   8'd106;
	gem_pad_to_csc_hs_me1b_odd[ 29]     =   8'd105;
	gem_pad_to_csc_hs_me1b_odd[ 30]     =   8'd105;
	gem_pad_to_csc_hs_me1b_odd[ 31]     =   8'd104;
	gem_pad_to_csc_hs_me1b_odd[ 32]     =   8'd103;
	gem_pad_to_csc_hs_me1b_odd[ 33]     =   8'd103;
	gem_pad_to_csc_hs_me1b_odd[ 34]     =   8'd102;
	gem_pad_to_csc_hs_me1b_odd[ 35]     =   8'd101;
	gem_pad_to_csc_hs_me1b_odd[ 36]     =   8'd101;
	gem_pad_to_csc_hs_me1b_odd[ 37]     =   8'd100;
	gem_pad_to_csc_hs_me1b_odd[ 38]     =   8'd100;
	gem_pad_to_csc_hs_me1b_odd[ 39]     =   8'd99;
	gem_pad_to_csc_hs_me1b_odd[ 40]     =   8'd98;
	gem_pad_to_csc_hs_me1b_odd[ 41]     =   8'd98;
	gem_pad_to_csc_hs_me1b_odd[ 42]     =   8'd97;
	gem_pad_to_csc_hs_me1b_odd[ 43]     =   8'd96;
	gem_pad_to_csc_hs_me1b_odd[ 44]     =   8'd96;
	gem_pad_to_csc_hs_me1b_odd[ 45]     =   8'd95;
	gem_pad_to_csc_hs_me1b_odd[ 46]     =   8'd95;
	gem_pad_to_csc_hs_me1b_odd[ 47]     =   8'd94;
	gem_pad_to_csc_hs_me1b_odd[ 48]     =   8'd93;
	gem_pad_to_csc_hs_me1b_odd[ 49]     =   8'd93;
	gem_pad_to_csc_hs_me1b_odd[ 50]     =   8'd92;
	gem_pad_to_csc_hs_me1b_odd[ 51]     =   8'd91;
	gem_pad_to_csc_hs_me1b_odd[ 52]     =   8'd91;
	gem_pad_to_csc_hs_me1b_odd[ 53]     =   8'd90;
	gem_pad_to_csc_hs_me1b_odd[ 54]     =   8'd90;
	gem_pad_to_csc_hs_me1b_odd[ 55]     =   8'd89;
	gem_pad_to_csc_hs_me1b_odd[ 56]     =   8'd88;
	gem_pad_to_csc_hs_me1b_odd[ 57]     =   8'd88;
	gem_pad_to_csc_hs_me1b_odd[ 58]     =   8'd87;
	gem_pad_to_csc_hs_me1b_odd[ 59]     =   8'd86;
	gem_pad_to_csc_hs_me1b_odd[ 60]     =   8'd86;
	gem_pad_to_csc_hs_me1b_odd[ 61]     =   8'd85;
	gem_pad_to_csc_hs_me1b_odd[ 62]     =   8'd85;
	gem_pad_to_csc_hs_me1b_odd[ 63]     =   8'd84;
	gem_pad_to_csc_hs_me1b_odd[ 64]     =   8'd83;
	gem_pad_to_csc_hs_me1b_odd[ 65]     =   8'd83;
	gem_pad_to_csc_hs_me1b_odd[ 66]     =   8'd82;
	gem_pad_to_csc_hs_me1b_odd[ 67]     =   8'd81;
	gem_pad_to_csc_hs_me1b_odd[ 68]     =   8'd81;
	gem_pad_to_csc_hs_me1b_odd[ 69]     =   8'd80;
	gem_pad_to_csc_hs_me1b_odd[ 70]     =   8'd80;
	gem_pad_to_csc_hs_me1b_odd[ 71]     =   8'd79;
	gem_pad_to_csc_hs_me1b_odd[ 72]     =   8'd78;
	gem_pad_to_csc_hs_me1b_odd[ 73]     =   8'd78;
	gem_pad_to_csc_hs_me1b_odd[ 74]     =   8'd77;
	gem_pad_to_csc_hs_me1b_odd[ 75]     =   8'd76;
	gem_pad_to_csc_hs_me1b_odd[ 76]     =   8'd76;
	gem_pad_to_csc_hs_me1b_odd[ 77]     =   8'd75;
	gem_pad_to_csc_hs_me1b_odd[ 78]     =   8'd75;
	gem_pad_to_csc_hs_me1b_odd[ 79]     =   8'd74;
	gem_pad_to_csc_hs_me1b_odd[ 80]     =   8'd73;
	gem_pad_to_csc_hs_me1b_odd[ 81]     =   8'd73;
	gem_pad_to_csc_hs_me1b_odd[ 82]     =   8'd72;
	gem_pad_to_csc_hs_me1b_odd[ 83]     =   8'd71;
	gem_pad_to_csc_hs_me1b_odd[ 84]     =   8'd71;
	gem_pad_to_csc_hs_me1b_odd[ 85]     =   8'd70;
	gem_pad_to_csc_hs_me1b_odd[ 86]     =   8'd70;
	gem_pad_to_csc_hs_me1b_odd[ 87]     =   8'd69;
	gem_pad_to_csc_hs_me1b_odd[ 88]     =   8'd68;
	gem_pad_to_csc_hs_me1b_odd[ 89]     =   8'd68;
	gem_pad_to_csc_hs_me1b_odd[ 90]     =   8'd67;
	gem_pad_to_csc_hs_me1b_odd[ 91]     =   8'd66;
	gem_pad_to_csc_hs_me1b_odd[ 92]     =   8'd66;
	gem_pad_to_csc_hs_me1b_odd[ 93]     =   8'd65;
	gem_pad_to_csc_hs_me1b_odd[ 94]     =   8'd65;
	gem_pad_to_csc_hs_me1b_odd[ 95]     =   8'd64;
	gem_pad_to_csc_hs_me1b_odd[ 96]     =   8'd63;
	gem_pad_to_csc_hs_me1b_odd[ 97]     =   8'd63;
	gem_pad_to_csc_hs_me1b_odd[ 98]     =   8'd62;
	gem_pad_to_csc_hs_me1b_odd[ 99]     =   8'd61;
	gem_pad_to_csc_hs_me1b_odd[100]     =   8'd61;
	gem_pad_to_csc_hs_me1b_odd[101]     =   8'd60;
	gem_pad_to_csc_hs_me1b_odd[102]     =   8'd60;
	gem_pad_to_csc_hs_me1b_odd[103]     =   8'd59;
	gem_pad_to_csc_hs_me1b_odd[104]     =   8'd58;
	gem_pad_to_csc_hs_me1b_odd[105]     =   8'd58;
	gem_pad_to_csc_hs_me1b_odd[106]     =   8'd57;
	gem_pad_to_csc_hs_me1b_odd[107]     =   8'd56;
	gem_pad_to_csc_hs_me1b_odd[108]     =   8'd56;
	gem_pad_to_csc_hs_me1b_odd[109]     =   8'd55;
	gem_pad_to_csc_hs_me1b_odd[110]     =   8'd55;
	gem_pad_to_csc_hs_me1b_odd[111]     =   8'd54;
	gem_pad_to_csc_hs_me1b_odd[112]     =   8'd53;
	gem_pad_to_csc_hs_me1b_odd[113]     =   8'd53;
	gem_pad_to_csc_hs_me1b_odd[114]     =   8'd52;
	gem_pad_to_csc_hs_me1b_odd[115]     =   8'd51;
	gem_pad_to_csc_hs_me1b_odd[116]     =   8'd51;
	gem_pad_to_csc_hs_me1b_odd[117]     =   8'd50;
	gem_pad_to_csc_hs_me1b_odd[118]     =   8'd50;
	gem_pad_to_csc_hs_me1b_odd[119]     =   8'd49;
	gem_pad_to_csc_hs_me1b_odd[120]     =   8'd48;
	gem_pad_to_csc_hs_me1b_odd[121]     =   8'd48;
	gem_pad_to_csc_hs_me1b_odd[122]     =   8'd47;
	gem_pad_to_csc_hs_me1b_odd[123]     =   8'd46;
	gem_pad_to_csc_hs_me1b_odd[124]     =   8'd46;
	gem_pad_to_csc_hs_me1b_odd[125]     =   8'd45;
	gem_pad_to_csc_hs_me1b_odd[126]     =   8'd45;
	gem_pad_to_csc_hs_me1b_odd[127]     =   8'd44;
	gem_pad_to_csc_hs_me1b_odd[128]     =   8'd43;
	gem_pad_to_csc_hs_me1b_odd[129]     =   8'd43;
	gem_pad_to_csc_hs_me1b_odd[130]     =   8'd42;
	gem_pad_to_csc_hs_me1b_odd[131]     =   8'd41;
	gem_pad_to_csc_hs_me1b_odd[132]     =   8'd41;
	gem_pad_to_csc_hs_me1b_odd[133]     =   8'd40;
	gem_pad_to_csc_hs_me1b_odd[134]     =   8'd40;
	gem_pad_to_csc_hs_me1b_odd[135]     =   8'd39;
	gem_pad_to_csc_hs_me1b_odd[136]     =   8'd38;
	gem_pad_to_csc_hs_me1b_odd[137]     =   8'd38;
	gem_pad_to_csc_hs_me1b_odd[138]     =   8'd37;
	gem_pad_to_csc_hs_me1b_odd[139]     =   8'd36;
	gem_pad_to_csc_hs_me1b_odd[140]     =   8'd36;
	gem_pad_to_csc_hs_me1b_odd[141]     =   8'd35;
	gem_pad_to_csc_hs_me1b_odd[142]     =   8'd35;
	gem_pad_to_csc_hs_me1b_odd[143]     =   8'd34;
	gem_pad_to_csc_hs_me1b_odd[144]     =   8'd33;
	gem_pad_to_csc_hs_me1b_odd[145]     =   8'd33;
	gem_pad_to_csc_hs_me1b_odd[146]     =   8'd32;
	gem_pad_to_csc_hs_me1b_odd[147]     =   8'd31;
	gem_pad_to_csc_hs_me1b_odd[148]     =   8'd31;
	gem_pad_to_csc_hs_me1b_odd[149]     =   8'd30;
	gem_pad_to_csc_hs_me1b_odd[150]     =   8'd30;
	gem_pad_to_csc_hs_me1b_odd[151]     =   8'd29;
	gem_pad_to_csc_hs_me1b_odd[152]     =   8'd28;
	gem_pad_to_csc_hs_me1b_odd[153]     =   8'd28;
	gem_pad_to_csc_hs_me1b_odd[154]     =   8'd27;
	gem_pad_to_csc_hs_me1b_odd[155]     =   8'd26;
	gem_pad_to_csc_hs_me1b_odd[156]     =   8'd26;
	gem_pad_to_csc_hs_me1b_odd[157]     =   8'd25;
	gem_pad_to_csc_hs_me1b_odd[158]     =   8'd25;
	gem_pad_to_csc_hs_me1b_odd[159]     =   8'd24;
	gem_pad_to_csc_hs_me1b_odd[160]     =   8'd23;
	gem_pad_to_csc_hs_me1b_odd[161]     =   8'd23;
	gem_pad_to_csc_hs_me1b_odd[162]     =   8'd22;
	gem_pad_to_csc_hs_me1b_odd[163]     =   8'd21;
	gem_pad_to_csc_hs_me1b_odd[164]     =   8'd21;
	gem_pad_to_csc_hs_me1b_odd[165]     =   8'd20;
	gem_pad_to_csc_hs_me1b_odd[166]     =   8'd20;
	gem_pad_to_csc_hs_me1b_odd[167]     =   8'd19;
	gem_pad_to_csc_hs_me1b_odd[168]     =   8'd18;
	gem_pad_to_csc_hs_me1b_odd[169]     =   8'd18;
	gem_pad_to_csc_hs_me1b_odd[170]     =   8'd17;
	gem_pad_to_csc_hs_me1b_odd[171]     =   8'd16;
	gem_pad_to_csc_hs_me1b_odd[172]     =   8'd16;
	gem_pad_to_csc_hs_me1b_odd[173]     =   8'd15;
	gem_pad_to_csc_hs_me1b_odd[174]     =   8'd15;
	gem_pad_to_csc_hs_me1b_odd[175]     =   8'd14;
	gem_pad_to_csc_hs_me1b_odd[176]     =   8'd13;
	gem_pad_to_csc_hs_me1b_odd[177]     =   8'd13;
	gem_pad_to_csc_hs_me1b_odd[178]     =   8'd12;
	gem_pad_to_csc_hs_me1b_odd[179]     =   8'd11;
	gem_pad_to_csc_hs_me1b_odd[180]     =   8'd11;
	gem_pad_to_csc_hs_me1b_odd[181]     =   8'd10;
	gem_pad_to_csc_hs_me1b_odd[182]     =   8'd10;
	gem_pad_to_csc_hs_me1b_odd[183]     =   8'd9;
	gem_pad_to_csc_hs_me1b_odd[184]     =   8'd8;
	gem_pad_to_csc_hs_me1b_odd[185]     =   8'd8;
	gem_pad_to_csc_hs_me1b_odd[186]     =   8'd7;
	gem_pad_to_csc_hs_me1b_odd[187]     =   8'd7;
	gem_pad_to_csc_hs_me1b_odd[188]     =   8'd6;
	gem_pad_to_csc_hs_me1b_odd[189]     =   8'd5;
	gem_pad_to_csc_hs_me1b_odd[190]     =   8'd5;
	gem_pad_to_csc_hs_me1b_odd[191]     =   8'd4;
  end


  initial begin
	gem_pad_to_csc_hs_me1b_even[  0]     =   8'd4;
	gem_pad_to_csc_hs_me1b_even[  1]     =   8'd4;
	gem_pad_to_csc_hs_me1b_even[  2]     =   8'd5;
	gem_pad_to_csc_hs_me1b_even[  3]     =   8'd6;
	gem_pad_to_csc_hs_me1b_even[  4]     =   8'd6;
	gem_pad_to_csc_hs_me1b_even[  5]     =   8'd7;
	gem_pad_to_csc_hs_me1b_even[  6]     =   8'd7;
	gem_pad_to_csc_hs_me1b_even[  7]     =   8'd8;
	gem_pad_to_csc_hs_me1b_even[  8]     =   8'd9;
	gem_pad_to_csc_hs_me1b_even[  9]     =   8'd9;
	gem_pad_to_csc_hs_me1b_even[ 10]     =   8'd10;
	gem_pad_to_csc_hs_me1b_even[ 11]     =   8'd11;
	gem_pad_to_csc_hs_me1b_even[ 12]     =   8'd11;
	gem_pad_to_csc_hs_me1b_even[ 13]     =   8'd12;
	gem_pad_to_csc_hs_me1b_even[ 14]     =   8'd12;
	gem_pad_to_csc_hs_me1b_even[ 15]     =   8'd13;
	gem_pad_to_csc_hs_me1b_even[ 16]     =   8'd14;
	gem_pad_to_csc_hs_me1b_even[ 17]     =   8'd14;
	gem_pad_to_csc_hs_me1b_even[ 18]     =   8'd15;
	gem_pad_to_csc_hs_me1b_even[ 19]     =   8'd16;
	gem_pad_to_csc_hs_me1b_even[ 20]     =   8'd16;
	gem_pad_to_csc_hs_me1b_even[ 21]     =   8'd17;
	gem_pad_to_csc_hs_me1b_even[ 22]     =   8'd17;
	gem_pad_to_csc_hs_me1b_even[ 23]     =   8'd18;
	gem_pad_to_csc_hs_me1b_even[ 24]     =   8'd19;
	gem_pad_to_csc_hs_me1b_even[ 25]     =   8'd19;
	gem_pad_to_csc_hs_me1b_even[ 26]     =   8'd20;
	gem_pad_to_csc_hs_me1b_even[ 27]     =   8'd20;
	gem_pad_to_csc_hs_me1b_even[ 28]     =   8'd21;
	gem_pad_to_csc_hs_me1b_even[ 29]     =   8'd22;
	gem_pad_to_csc_hs_me1b_even[ 30]     =   8'd22;
	gem_pad_to_csc_hs_me1b_even[ 31]     =   8'd23;
	gem_pad_to_csc_hs_me1b_even[ 32]     =   8'd24;
	gem_pad_to_csc_hs_me1b_even[ 33]     =   8'd24;
	gem_pad_to_csc_hs_me1b_even[ 34]     =   8'd25;
	gem_pad_to_csc_hs_me1b_even[ 35]     =   8'd25;
	gem_pad_to_csc_hs_me1b_even[ 36]     =   8'd26;
	gem_pad_to_csc_hs_me1b_even[ 37]     =   8'd27;
	gem_pad_to_csc_hs_me1b_even[ 38]     =   8'd27;
	gem_pad_to_csc_hs_me1b_even[ 39]     =   8'd28;
	gem_pad_to_csc_hs_me1b_even[ 40]     =   8'd29;
	gem_pad_to_csc_hs_me1b_even[ 41]     =   8'd29;
	gem_pad_to_csc_hs_me1b_even[ 42]     =   8'd30;
	gem_pad_to_csc_hs_me1b_even[ 43]     =   8'd30;
	gem_pad_to_csc_hs_me1b_even[ 44]     =   8'd31;
	gem_pad_to_csc_hs_me1b_even[ 45]     =   8'd32;
	gem_pad_to_csc_hs_me1b_even[ 46]     =   8'd32;
	gem_pad_to_csc_hs_me1b_even[ 47]     =   8'd33;
	gem_pad_to_csc_hs_me1b_even[ 48]     =   8'd34;
	gem_pad_to_csc_hs_me1b_even[ 49]     =   8'd34;
	gem_pad_to_csc_hs_me1b_even[ 50]     =   8'd35;
	gem_pad_to_csc_hs_me1b_even[ 51]     =   8'd35;
	gem_pad_to_csc_hs_me1b_even[ 52]     =   8'd36;
	gem_pad_to_csc_hs_me1b_even[ 53]     =   8'd37;
	gem_pad_to_csc_hs_me1b_even[ 54]     =   8'd37;
	gem_pad_to_csc_hs_me1b_even[ 55]     =   8'd38;
	gem_pad_to_csc_hs_me1b_even[ 56]     =   8'd39;
	gem_pad_to_csc_hs_me1b_even[ 57]     =   8'd39;
	gem_pad_to_csc_hs_me1b_even[ 58]     =   8'd40;
	gem_pad_to_csc_hs_me1b_even[ 59]     =   8'd40;
	gem_pad_to_csc_hs_me1b_even[ 60]     =   8'd41;
	gem_pad_to_csc_hs_me1b_even[ 61]     =   8'd42;
	gem_pad_to_csc_hs_me1b_even[ 62]     =   8'd42;
	gem_pad_to_csc_hs_me1b_even[ 63]     =   8'd43;
	gem_pad_to_csc_hs_me1b_even[ 64]     =   8'd44;
	gem_pad_to_csc_hs_me1b_even[ 65]     =   8'd44;
	gem_pad_to_csc_hs_me1b_even[ 66]     =   8'd45;
	gem_pad_to_csc_hs_me1b_even[ 67]     =   8'd45;
	gem_pad_to_csc_hs_me1b_even[ 68]     =   8'd46;
	gem_pad_to_csc_hs_me1b_even[ 69]     =   8'd47;
	gem_pad_to_csc_hs_me1b_even[ 70]     =   8'd47;
	gem_pad_to_csc_hs_me1b_even[ 71]     =   8'd48;
	gem_pad_to_csc_hs_me1b_even[ 72]     =   8'd49;
	gem_pad_to_csc_hs_me1b_even[ 73]     =   8'd49;
	gem_pad_to_csc_hs_me1b_even[ 74]     =   8'd50;
	gem_pad_to_csc_hs_me1b_even[ 75]     =   8'd50;
	gem_pad_to_csc_hs_me1b_even[ 76]     =   8'd51;
	gem_pad_to_csc_hs_me1b_even[ 77]     =   8'd52;
	gem_pad_to_csc_hs_me1b_even[ 78]     =   8'd52;
	gem_pad_to_csc_hs_me1b_even[ 79]     =   8'd53;
	gem_pad_to_csc_hs_me1b_even[ 80]     =   8'd54;
	gem_pad_to_csc_hs_me1b_even[ 81]     =   8'd54;
	gem_pad_to_csc_hs_me1b_even[ 82]     =   8'd55;
	gem_pad_to_csc_hs_me1b_even[ 83]     =   8'd55;
	gem_pad_to_csc_hs_me1b_even[ 84]     =   8'd56;
	gem_pad_to_csc_hs_me1b_even[ 85]     =   8'd57;
	gem_pad_to_csc_hs_me1b_even[ 86]     =   8'd57;
	gem_pad_to_csc_hs_me1b_even[ 87]     =   8'd58;
	gem_pad_to_csc_hs_me1b_even[ 88]     =   8'd59;
	gem_pad_to_csc_hs_me1b_even[ 89]     =   8'd59;
	gem_pad_to_csc_hs_me1b_even[ 90]     =   8'd60;
	gem_pad_to_csc_hs_me1b_even[ 91]     =   8'd60;
	gem_pad_to_csc_hs_me1b_even[ 92]     =   8'd61;
	gem_pad_to_csc_hs_me1b_even[ 93]     =   8'd62;
	gem_pad_to_csc_hs_me1b_even[ 94]     =   8'd62;
	gem_pad_to_csc_hs_me1b_even[ 95]     =   8'd63;
	gem_pad_to_csc_hs_me1b_even[ 96]     =   8'd64;
	gem_pad_to_csc_hs_me1b_even[ 97]     =   8'd64;
	gem_pad_to_csc_hs_me1b_even[ 98]     =   8'd65;
	gem_pad_to_csc_hs_me1b_even[ 99]     =   8'd65;
	gem_pad_to_csc_hs_me1b_even[100]     =   8'd66;
	gem_pad_to_csc_hs_me1b_even[101]     =   8'd67;
	gem_pad_to_csc_hs_me1b_even[102]     =   8'd67;
	gem_pad_to_csc_hs_me1b_even[103]     =   8'd68;
	gem_pad_to_csc_hs_me1b_even[104]     =   8'd69;
	gem_pad_to_csc_hs_me1b_even[105]     =   8'd69;
	gem_pad_to_csc_hs_me1b_even[106]     =   8'd70;
	gem_pad_to_csc_hs_me1b_even[107]     =   8'd70;
	gem_pad_to_csc_hs_me1b_even[108]     =   8'd71;
	gem_pad_to_csc_hs_me1b_even[109]     =   8'd72;
	gem_pad_to_csc_hs_me1b_even[110]     =   8'd72;
	gem_pad_to_csc_hs_me1b_even[111]     =   8'd73;
	gem_pad_to_csc_hs_me1b_even[112]     =   8'd74;
	gem_pad_to_csc_hs_me1b_even[113]     =   8'd74;
	gem_pad_to_csc_hs_me1b_even[114]     =   8'd75;
	gem_pad_to_csc_hs_me1b_even[115]     =   8'd75;
	gem_pad_to_csc_hs_me1b_even[116]     =   8'd76;
	gem_pad_to_csc_hs_me1b_even[117]     =   8'd77;
	gem_pad_to_csc_hs_me1b_even[118]     =   8'd77;
	gem_pad_to_csc_hs_me1b_even[119]     =   8'd78;
	gem_pad_to_csc_hs_me1b_even[120]     =   8'd79;
	gem_pad_to_csc_hs_me1b_even[121]     =   8'd79;
	gem_pad_to_csc_hs_me1b_even[122]     =   8'd80;
	gem_pad_to_csc_hs_me1b_even[123]     =   8'd80;
	gem_pad_to_csc_hs_me1b_even[124]     =   8'd81;
	gem_pad_to_csc_hs_me1b_even[125]     =   8'd82;
	gem_pad_to_csc_hs_me1b_even[126]     =   8'd82;
	gem_pad_to_csc_hs_me1b_even[127]     =   8'd83;
	gem_pad_to_csc_hs_me1b_even[128]     =   8'd84;
	gem_pad_to_csc_hs_me1b_even[129]     =   8'd84;
	gem_pad_to_csc_hs_me1b_even[130]     =   8'd85;
	gem_pad_to_csc_hs_me1b_even[131]     =   8'd85;
	gem_pad_to_csc_hs_me1b_even[132]     =   8'd86;
	gem_pad_to_csc_hs_me1b_even[133]     =   8'd87;
	gem_pad_to_csc_hs_me1b_even[134]     =   8'd87;
	gem_pad_to_csc_hs_me1b_even[135]     =   8'd88;
	gem_pad_to_csc_hs_me1b_even[136]     =   8'd89;
	gem_pad_to_csc_hs_me1b_even[137]     =   8'd89;
	gem_pad_to_csc_hs_me1b_even[138]     =   8'd90;
	gem_pad_to_csc_hs_me1b_even[139]     =   8'd90;
	gem_pad_to_csc_hs_me1b_even[140]     =   8'd91;
	gem_pad_to_csc_hs_me1b_even[141]     =   8'd92;
	gem_pad_to_csc_hs_me1b_even[142]     =   8'd92;
	gem_pad_to_csc_hs_me1b_even[143]     =   8'd93;
	gem_pad_to_csc_hs_me1b_even[144]     =   8'd94;
	gem_pad_to_csc_hs_me1b_even[145]     =   8'd94;
	gem_pad_to_csc_hs_me1b_even[146]     =   8'd95;
	gem_pad_to_csc_hs_me1b_even[147]     =   8'd95;
	gem_pad_to_csc_hs_me1b_even[148]     =   8'd96;
	gem_pad_to_csc_hs_me1b_even[149]     =   8'd97;
	gem_pad_to_csc_hs_me1b_even[150]     =   8'd97;
	gem_pad_to_csc_hs_me1b_even[151]     =   8'd98;
	gem_pad_to_csc_hs_me1b_even[152]     =   8'd99;
	gem_pad_to_csc_hs_me1b_even[153]     =   8'd99;
	gem_pad_to_csc_hs_me1b_even[154]     =   8'd100;
	gem_pad_to_csc_hs_me1b_even[155]     =   8'd100;
	gem_pad_to_csc_hs_me1b_even[156]     =   8'd101;
	gem_pad_to_csc_hs_me1b_even[157]     =   8'd102;
	gem_pad_to_csc_hs_me1b_even[158]     =   8'd102;
	gem_pad_to_csc_hs_me1b_even[159]     =   8'd103;
	gem_pad_to_csc_hs_me1b_even[160]     =   8'd104;
	gem_pad_to_csc_hs_me1b_even[161]     =   8'd104;
	gem_pad_to_csc_hs_me1b_even[162]     =   8'd105;
	gem_pad_to_csc_hs_me1b_even[163]     =   8'd105;
	gem_pad_to_csc_hs_me1b_even[164]     =   8'd106;
	gem_pad_to_csc_hs_me1b_even[165]     =   8'd107;
	gem_pad_to_csc_hs_me1b_even[166]     =   8'd107;
	gem_pad_to_csc_hs_me1b_even[167]     =   8'd108;
	gem_pad_to_csc_hs_me1b_even[168]     =   8'd109;
	gem_pad_to_csc_hs_me1b_even[169]     =   8'd109;
	gem_pad_to_csc_hs_me1b_even[170]     =   8'd110;
	gem_pad_to_csc_hs_me1b_even[171]     =   8'd110;
	gem_pad_to_csc_hs_me1b_even[172]     =   8'd111;
	gem_pad_to_csc_hs_me1b_even[173]     =   8'd112;
	gem_pad_to_csc_hs_me1b_even[174]     =   8'd112;
	gem_pad_to_csc_hs_me1b_even[175]     =   8'd113;
	gem_pad_to_csc_hs_me1b_even[176]     =   8'd114;
	gem_pad_to_csc_hs_me1b_even[177]     =   8'd114;
	gem_pad_to_csc_hs_me1b_even[178]     =   8'd115;
	gem_pad_to_csc_hs_me1b_even[179]     =   8'd115;
	gem_pad_to_csc_hs_me1b_even[180]     =   8'd116;
	gem_pad_to_csc_hs_me1b_even[181]     =   8'd117;
	gem_pad_to_csc_hs_me1b_even[182]     =   8'd117;
	gem_pad_to_csc_hs_me1b_even[183]     =   8'd118;
	gem_pad_to_csc_hs_me1b_even[184]     =   8'd119;
	gem_pad_to_csc_hs_me1b_even[185]     =   8'd119;
	gem_pad_to_csc_hs_me1b_even[186]     =   8'd120;
	gem_pad_to_csc_hs_me1b_even[187]     =   8'd120;
	gem_pad_to_csc_hs_me1b_even[188]     =   8'd121;
	gem_pad_to_csc_hs_me1b_even[189]     =   8'd122;
	gem_pad_to_csc_hs_me1b_even[190]     =   8'd122;
	gem_pad_to_csc_hs_me1b_even[191]     =   8'd123;
  end


  initial begin
	gem_pad_to_csc_hs_me1a_odd[  0]     =   8'd221;
	gem_pad_to_csc_hs_me1a_odd[  1]     =   8'd220;
	gem_pad_to_csc_hs_me1a_odd[  2]     =   8'd220;
	gem_pad_to_csc_hs_me1a_odd[  3]     =   8'd220;
	gem_pad_to_csc_hs_me1a_odd[  4]     =   8'd219;
	gem_pad_to_csc_hs_me1a_odd[  5]     =   8'd219;
	gem_pad_to_csc_hs_me1a_odd[  6]     =   8'd218;
	gem_pad_to_csc_hs_me1a_odd[  7]     =   8'd218;
	gem_pad_to_csc_hs_me1a_odd[  8]     =   8'd217;
	gem_pad_to_csc_hs_me1a_odd[  9]     =   8'd217;
	gem_pad_to_csc_hs_me1a_odd[ 10]     =   8'd216;
	gem_pad_to_csc_hs_me1a_odd[ 11]     =   8'd216;
	gem_pad_to_csc_hs_me1a_odd[ 12]     =   8'd215;
	gem_pad_to_csc_hs_me1a_odd[ 13]     =   8'd215;
	gem_pad_to_csc_hs_me1a_odd[ 14]     =   8'd214;
	gem_pad_to_csc_hs_me1a_odd[ 15]     =   8'd214;
	gem_pad_to_csc_hs_me1a_odd[ 16]     =   8'd213;
	gem_pad_to_csc_hs_me1a_odd[ 17]     =   8'd213;
	gem_pad_to_csc_hs_me1a_odd[ 18]     =   8'd212;
	gem_pad_to_csc_hs_me1a_odd[ 19]     =   8'd212;
	gem_pad_to_csc_hs_me1a_odd[ 20]     =   8'd211;
	gem_pad_to_csc_hs_me1a_odd[ 21]     =   8'd211;
	gem_pad_to_csc_hs_me1a_odd[ 22]     =   8'd211;
	gem_pad_to_csc_hs_me1a_odd[ 23]     =   8'd210;
	gem_pad_to_csc_hs_me1a_odd[ 24]     =   8'd210;
	gem_pad_to_csc_hs_me1a_odd[ 25]     =   8'd209;
	gem_pad_to_csc_hs_me1a_odd[ 26]     =   8'd209;
	gem_pad_to_csc_hs_me1a_odd[ 27]     =   8'd208;
	gem_pad_to_csc_hs_me1a_odd[ 28]     =   8'd208;
	gem_pad_to_csc_hs_me1a_odd[ 29]     =   8'd207;
	gem_pad_to_csc_hs_me1a_odd[ 30]     =   8'd207;
	gem_pad_to_csc_hs_me1a_odd[ 31]     =   8'd206;
	gem_pad_to_csc_hs_me1a_odd[ 32]     =   8'd206;
	gem_pad_to_csc_hs_me1a_odd[ 33]     =   8'd205;
	gem_pad_to_csc_hs_me1a_odd[ 34]     =   8'd205;
	gem_pad_to_csc_hs_me1a_odd[ 35]     =   8'd204;
	gem_pad_to_csc_hs_me1a_odd[ 36]     =   8'd204;
	gem_pad_to_csc_hs_me1a_odd[ 37]     =   8'd203;
	gem_pad_to_csc_hs_me1a_odd[ 38]     =   8'd203;
	gem_pad_to_csc_hs_me1a_odd[ 39]     =   8'd202;
	gem_pad_to_csc_hs_me1a_odd[ 40]     =   8'd202;
	gem_pad_to_csc_hs_me1a_odd[ 41]     =   8'd201;
	gem_pad_to_csc_hs_me1a_odd[ 42]     =   8'd201;
	gem_pad_to_csc_hs_me1a_odd[ 43]     =   8'd201;
	gem_pad_to_csc_hs_me1a_odd[ 44]     =   8'd200;
	gem_pad_to_csc_hs_me1a_odd[ 45]     =   8'd200;
	gem_pad_to_csc_hs_me1a_odd[ 46]     =   8'd199;
	gem_pad_to_csc_hs_me1a_odd[ 47]     =   8'd199;
	gem_pad_to_csc_hs_me1a_odd[ 48]     =   8'd198;
	gem_pad_to_csc_hs_me1a_odd[ 49]     =   8'd198;
	gem_pad_to_csc_hs_me1a_odd[ 50]     =   8'd197;
	gem_pad_to_csc_hs_me1a_odd[ 51]     =   8'd197;
	gem_pad_to_csc_hs_me1a_odd[ 52]     =   8'd196;
	gem_pad_to_csc_hs_me1a_odd[ 53]     =   8'd196;
	gem_pad_to_csc_hs_me1a_odd[ 54]     =   8'd195;
	gem_pad_to_csc_hs_me1a_odd[ 55]     =   8'd195;
	gem_pad_to_csc_hs_me1a_odd[ 56]     =   8'd194;
	gem_pad_to_csc_hs_me1a_odd[ 57]     =   8'd194;
	gem_pad_to_csc_hs_me1a_odd[ 58]     =   8'd193;
	gem_pad_to_csc_hs_me1a_odd[ 59]     =   8'd193;
	gem_pad_to_csc_hs_me1a_odd[ 60]     =   8'd192;
	gem_pad_to_csc_hs_me1a_odd[ 61]     =   8'd192;
	gem_pad_to_csc_hs_me1a_odd[ 62]     =   8'd191;
	gem_pad_to_csc_hs_me1a_odd[ 63]     =   8'd191;
	gem_pad_to_csc_hs_me1a_odd[ 64]     =   8'd191;
	gem_pad_to_csc_hs_me1a_odd[ 65]     =   8'd190;
	gem_pad_to_csc_hs_me1a_odd[ 66]     =   8'd190;
	gem_pad_to_csc_hs_me1a_odd[ 67]     =   8'd189;
	gem_pad_to_csc_hs_me1a_odd[ 68]     =   8'd189;
	gem_pad_to_csc_hs_me1a_odd[ 69]     =   8'd188;
	gem_pad_to_csc_hs_me1a_odd[ 70]     =   8'd188;
	gem_pad_to_csc_hs_me1a_odd[ 71]     =   8'd187;
	gem_pad_to_csc_hs_me1a_odd[ 72]     =   8'd187;
	gem_pad_to_csc_hs_me1a_odd[ 73]     =   8'd186;
	gem_pad_to_csc_hs_me1a_odd[ 74]     =   8'd186;
	gem_pad_to_csc_hs_me1a_odd[ 75]     =   8'd185;
	gem_pad_to_csc_hs_me1a_odd[ 76]     =   8'd185;
	gem_pad_to_csc_hs_me1a_odd[ 77]     =   8'd184;
	gem_pad_to_csc_hs_me1a_odd[ 78]     =   8'd184;
	gem_pad_to_csc_hs_me1a_odd[ 79]     =   8'd183;
	gem_pad_to_csc_hs_me1a_odd[ 80]     =   8'd183;
	gem_pad_to_csc_hs_me1a_odd[ 81]     =   8'd182;
	gem_pad_to_csc_hs_me1a_odd[ 82]     =   8'd182;
	gem_pad_to_csc_hs_me1a_odd[ 83]     =   8'd181;
	gem_pad_to_csc_hs_me1a_odd[ 84]     =   8'd181;
	gem_pad_to_csc_hs_me1a_odd[ 85]     =   8'd181;
	gem_pad_to_csc_hs_me1a_odd[ 86]     =   8'd180;
	gem_pad_to_csc_hs_me1a_odd[ 87]     =   8'd180;
	gem_pad_to_csc_hs_me1a_odd[ 88]     =   8'd179;
	gem_pad_to_csc_hs_me1a_odd[ 89]     =   8'd179;
	gem_pad_to_csc_hs_me1a_odd[ 90]     =   8'd178;
	gem_pad_to_csc_hs_me1a_odd[ 91]     =   8'd178;
	gem_pad_to_csc_hs_me1a_odd[ 92]     =   8'd177;
	gem_pad_to_csc_hs_me1a_odd[ 93]     =   8'd177;
	gem_pad_to_csc_hs_me1a_odd[ 94]     =   8'd176;
	gem_pad_to_csc_hs_me1a_odd[ 95]     =   8'd176;
	gem_pad_to_csc_hs_me1a_odd[ 96]     =   8'd175;
	gem_pad_to_csc_hs_me1a_odd[ 97]     =   8'd175;
	gem_pad_to_csc_hs_me1a_odd[ 98]     =   8'd174;
	gem_pad_to_csc_hs_me1a_odd[ 99]     =   8'd174;
	gem_pad_to_csc_hs_me1a_odd[100]     =   8'd173;
	gem_pad_to_csc_hs_me1a_odd[101]     =   8'd173;
	gem_pad_to_csc_hs_me1a_odd[102]     =   8'd172;
	gem_pad_to_csc_hs_me1a_odd[103]     =   8'd172;
	gem_pad_to_csc_hs_me1a_odd[104]     =   8'd171;
	gem_pad_to_csc_hs_me1a_odd[105]     =   8'd171;
	gem_pad_to_csc_hs_me1a_odd[106]     =   8'd171;
	gem_pad_to_csc_hs_me1a_odd[107]     =   8'd170;
	gem_pad_to_csc_hs_me1a_odd[108]     =   8'd170;
	gem_pad_to_csc_hs_me1a_odd[109]     =   8'd169;
	gem_pad_to_csc_hs_me1a_odd[110]     =   8'd169;
	gem_pad_to_csc_hs_me1a_odd[111]     =   8'd168;
	gem_pad_to_csc_hs_me1a_odd[112]     =   8'd168;
	gem_pad_to_csc_hs_me1a_odd[113]     =   8'd167;
	gem_pad_to_csc_hs_me1a_odd[114]     =   8'd167;
	gem_pad_to_csc_hs_me1a_odd[115]     =   8'd166;
	gem_pad_to_csc_hs_me1a_odd[116]     =   8'd166;
	gem_pad_to_csc_hs_me1a_odd[117]     =   8'd165;
	gem_pad_to_csc_hs_me1a_odd[118]     =   8'd165;
	gem_pad_to_csc_hs_me1a_odd[119]     =   8'd164;
	gem_pad_to_csc_hs_me1a_odd[120]     =   8'd164;
	gem_pad_to_csc_hs_me1a_odd[121]     =   8'd163;
	gem_pad_to_csc_hs_me1a_odd[122]     =   8'd163;
	gem_pad_to_csc_hs_me1a_odd[123]     =   8'd162;
	gem_pad_to_csc_hs_me1a_odd[124]     =   8'd162;
	gem_pad_to_csc_hs_me1a_odd[125]     =   8'd161;
	gem_pad_to_csc_hs_me1a_odd[126]     =   8'd161;
	gem_pad_to_csc_hs_me1a_odd[127]     =   8'd161;
	gem_pad_to_csc_hs_me1a_odd[128]     =   8'd160;
	gem_pad_to_csc_hs_me1a_odd[129]     =   8'd160;
	gem_pad_to_csc_hs_me1a_odd[130]     =   8'd159;
	gem_pad_to_csc_hs_me1a_odd[131]     =   8'd159;
	gem_pad_to_csc_hs_me1a_odd[132]     =   8'd158;
	gem_pad_to_csc_hs_me1a_odd[133]     =   8'd158;
	gem_pad_to_csc_hs_me1a_odd[134]     =   8'd157;
	gem_pad_to_csc_hs_me1a_odd[135]     =   8'd157;
	gem_pad_to_csc_hs_me1a_odd[136]     =   8'd156;
	gem_pad_to_csc_hs_me1a_odd[137]     =   8'd156;
	gem_pad_to_csc_hs_me1a_odd[138]     =   8'd155;
	gem_pad_to_csc_hs_me1a_odd[139]     =   8'd155;
	gem_pad_to_csc_hs_me1a_odd[140]     =   8'd154;
	gem_pad_to_csc_hs_me1a_odd[141]     =   8'd154;
	gem_pad_to_csc_hs_me1a_odd[142]     =   8'd153;
	gem_pad_to_csc_hs_me1a_odd[143]     =   8'd153;
	gem_pad_to_csc_hs_me1a_odd[144]     =   8'd152;
	gem_pad_to_csc_hs_me1a_odd[145]     =   8'd152;
	gem_pad_to_csc_hs_me1a_odd[146]     =   8'd151;
	gem_pad_to_csc_hs_me1a_odd[147]     =   8'd151;
	gem_pad_to_csc_hs_me1a_odd[148]     =   8'd151;
	gem_pad_to_csc_hs_me1a_odd[149]     =   8'd150;
	gem_pad_to_csc_hs_me1a_odd[150]     =   8'd150;
	gem_pad_to_csc_hs_me1a_odd[151]     =   8'd149;
	gem_pad_to_csc_hs_me1a_odd[152]     =   8'd149;
	gem_pad_to_csc_hs_me1a_odd[153]     =   8'd148;
	gem_pad_to_csc_hs_me1a_odd[154]     =   8'd148;
	gem_pad_to_csc_hs_me1a_odd[155]     =   8'd147;
	gem_pad_to_csc_hs_me1a_odd[156]     =   8'd147;
	gem_pad_to_csc_hs_me1a_odd[157]     =   8'd146;
	gem_pad_to_csc_hs_me1a_odd[158]     =   8'd146;
	gem_pad_to_csc_hs_me1a_odd[159]     =   8'd145;
	gem_pad_to_csc_hs_me1a_odd[160]     =   8'd145;
	gem_pad_to_csc_hs_me1a_odd[161]     =   8'd144;
	gem_pad_to_csc_hs_me1a_odd[162]     =   8'd144;
	gem_pad_to_csc_hs_me1a_odd[163]     =   8'd143;
	gem_pad_to_csc_hs_me1a_odd[164]     =   8'd143;
	gem_pad_to_csc_hs_me1a_odd[165]     =   8'd142;
	gem_pad_to_csc_hs_me1a_odd[166]     =   8'd142;
	gem_pad_to_csc_hs_me1a_odd[167]     =   8'd141;
	gem_pad_to_csc_hs_me1a_odd[168]     =   8'd141;
	gem_pad_to_csc_hs_me1a_odd[169]     =   8'd141;
	gem_pad_to_csc_hs_me1a_odd[170]     =   8'd140;
	gem_pad_to_csc_hs_me1a_odd[171]     =   8'd140;
	gem_pad_to_csc_hs_me1a_odd[172]     =   8'd139;
	gem_pad_to_csc_hs_me1a_odd[173]     =   8'd139;
	gem_pad_to_csc_hs_me1a_odd[174]     =   8'd138;
	gem_pad_to_csc_hs_me1a_odd[175]     =   8'd138;
	gem_pad_to_csc_hs_me1a_odd[176]     =   8'd137;
	gem_pad_to_csc_hs_me1a_odd[177]     =   8'd137;
	gem_pad_to_csc_hs_me1a_odd[178]     =   8'd136;
	gem_pad_to_csc_hs_me1a_odd[179]     =   8'd136;
	gem_pad_to_csc_hs_me1a_odd[180]     =   8'd135;
	gem_pad_to_csc_hs_me1a_odd[181]     =   8'd135;
	gem_pad_to_csc_hs_me1a_odd[182]     =   8'd134;
	gem_pad_to_csc_hs_me1a_odd[183]     =   8'd134;
	gem_pad_to_csc_hs_me1a_odd[184]     =   8'd133;
	gem_pad_to_csc_hs_me1a_odd[185]     =   8'd133;
	gem_pad_to_csc_hs_me1a_odd[186]     =   8'd132;
	gem_pad_to_csc_hs_me1a_odd[187]     =   8'd132;
	gem_pad_to_csc_hs_me1a_odd[188]     =   8'd132;
	gem_pad_to_csc_hs_me1a_odd[189]     =   8'd131;
	gem_pad_to_csc_hs_me1a_odd[190]     =   8'd131;
	gem_pad_to_csc_hs_me1a_odd[191]     =   8'd130;
  end

reg [ 7:0] gem_pad_to_csc_hs_me1a_even [191:0];

  initial begin
	gem_pad_to_csc_hs_me1a_even[  0]     =   8'd130;
	gem_pad_to_csc_hs_me1a_even[  1]     =   8'd131;
	gem_pad_to_csc_hs_me1a_even[  2]     =   8'd131;
	gem_pad_to_csc_hs_me1a_even[  3]     =   8'd131;
	gem_pad_to_csc_hs_me1a_even[  4]     =   8'd132;
	gem_pad_to_csc_hs_me1a_even[  5]     =   8'd132;
	gem_pad_to_csc_hs_me1a_even[  6]     =   8'd133;
	gem_pad_to_csc_hs_me1a_even[  7]     =   8'd133;
	gem_pad_to_csc_hs_me1a_even[  8]     =   8'd134;
	gem_pad_to_csc_hs_me1a_even[  9]     =   8'd134;
	gem_pad_to_csc_hs_me1a_even[ 10]     =   8'd135;
	gem_pad_to_csc_hs_me1a_even[ 11]     =   8'd135;
	gem_pad_to_csc_hs_me1a_even[ 12]     =   8'd136;
	gem_pad_to_csc_hs_me1a_even[ 13]     =   8'd136;
	gem_pad_to_csc_hs_me1a_even[ 14]     =   8'd137;
	gem_pad_to_csc_hs_me1a_even[ 15]     =   8'd137;
	gem_pad_to_csc_hs_me1a_even[ 16]     =   8'd138;
	gem_pad_to_csc_hs_me1a_even[ 17]     =   8'd138;
	gem_pad_to_csc_hs_me1a_even[ 18]     =   8'd139;
	gem_pad_to_csc_hs_me1a_even[ 19]     =   8'd139;
	gem_pad_to_csc_hs_me1a_even[ 20]     =   8'd140;
	gem_pad_to_csc_hs_me1a_even[ 21]     =   8'd140;
	gem_pad_to_csc_hs_me1a_even[ 22]     =   8'd140;
	gem_pad_to_csc_hs_me1a_even[ 23]     =   8'd141;
	gem_pad_to_csc_hs_me1a_even[ 24]     =   8'd141;
	gem_pad_to_csc_hs_me1a_even[ 25]     =   8'd142;
	gem_pad_to_csc_hs_me1a_even[ 26]     =   8'd142;
	gem_pad_to_csc_hs_me1a_even[ 27]     =   8'd143;
	gem_pad_to_csc_hs_me1a_even[ 28]     =   8'd143;
	gem_pad_to_csc_hs_me1a_even[ 29]     =   8'd144;
	gem_pad_to_csc_hs_me1a_even[ 30]     =   8'd144;
	gem_pad_to_csc_hs_me1a_even[ 31]     =   8'd145;
	gem_pad_to_csc_hs_me1a_even[ 32]     =   8'd145;
	gem_pad_to_csc_hs_me1a_even[ 33]     =   8'd146;
	gem_pad_to_csc_hs_me1a_even[ 34]     =   8'd146;
	gem_pad_to_csc_hs_me1a_even[ 35]     =   8'd147;
	gem_pad_to_csc_hs_me1a_even[ 36]     =   8'd147;
	gem_pad_to_csc_hs_me1a_even[ 37]     =   8'd148;
	gem_pad_to_csc_hs_me1a_even[ 38]     =   8'd148;
	gem_pad_to_csc_hs_me1a_even[ 39]     =   8'd149;
	gem_pad_to_csc_hs_me1a_even[ 40]     =   8'd149;
	gem_pad_to_csc_hs_me1a_even[ 41]     =   8'd150;
	gem_pad_to_csc_hs_me1a_even[ 42]     =   8'd150;
	gem_pad_to_csc_hs_me1a_even[ 43]     =   8'd150;
	gem_pad_to_csc_hs_me1a_even[ 44]     =   8'd151;
	gem_pad_to_csc_hs_me1a_even[ 45]     =   8'd151;
	gem_pad_to_csc_hs_me1a_even[ 46]     =   8'd152;
	gem_pad_to_csc_hs_me1a_even[ 47]     =   8'd152;
	gem_pad_to_csc_hs_me1a_even[ 48]     =   8'd153;
	gem_pad_to_csc_hs_me1a_even[ 49]     =   8'd153;
	gem_pad_to_csc_hs_me1a_even[ 50]     =   8'd154;
	gem_pad_to_csc_hs_me1a_even[ 51]     =   8'd154;
	gem_pad_to_csc_hs_me1a_even[ 52]     =   8'd155;
	gem_pad_to_csc_hs_me1a_even[ 53]     =   8'd155;
	gem_pad_to_csc_hs_me1a_even[ 54]     =   8'd156;
	gem_pad_to_csc_hs_me1a_even[ 55]     =   8'd156;
	gem_pad_to_csc_hs_me1a_even[ 56]     =   8'd157;
	gem_pad_to_csc_hs_me1a_even[ 57]     =   8'd157;
	gem_pad_to_csc_hs_me1a_even[ 58]     =   8'd158;
	gem_pad_to_csc_hs_me1a_even[ 59]     =   8'd158;
	gem_pad_to_csc_hs_me1a_even[ 60]     =   8'd159;
	gem_pad_to_csc_hs_me1a_even[ 61]     =   8'd159;
	gem_pad_to_csc_hs_me1a_even[ 62]     =   8'd160;
	gem_pad_to_csc_hs_me1a_even[ 63]     =   8'd160;
	gem_pad_to_csc_hs_me1a_even[ 64]     =   8'd160;
	gem_pad_to_csc_hs_me1a_even[ 65]     =   8'd161;
	gem_pad_to_csc_hs_me1a_even[ 66]     =   8'd161;
	gem_pad_to_csc_hs_me1a_even[ 67]     =   8'd162;
	gem_pad_to_csc_hs_me1a_even[ 68]     =   8'd162;
	gem_pad_to_csc_hs_me1a_even[ 69]     =   8'd163;
	gem_pad_to_csc_hs_me1a_even[ 70]     =   8'd163;
	gem_pad_to_csc_hs_me1a_even[ 71]     =   8'd164;
	gem_pad_to_csc_hs_me1a_even[ 72]     =   8'd164;
	gem_pad_to_csc_hs_me1a_even[ 73]     =   8'd165;
	gem_pad_to_csc_hs_me1a_even[ 74]     =   8'd165;
	gem_pad_to_csc_hs_me1a_even[ 75]     =   8'd166;
	gem_pad_to_csc_hs_me1a_even[ 76]     =   8'd166;
	gem_pad_to_csc_hs_me1a_even[ 77]     =   8'd167;
	gem_pad_to_csc_hs_me1a_even[ 78]     =   8'd167;
	gem_pad_to_csc_hs_me1a_even[ 79]     =   8'd168;
	gem_pad_to_csc_hs_me1a_even[ 80]     =   8'd168;
	gem_pad_to_csc_hs_me1a_even[ 81]     =   8'd169;
	gem_pad_to_csc_hs_me1a_even[ 82]     =   8'd169;
	gem_pad_to_csc_hs_me1a_even[ 83]     =   8'd170;
	gem_pad_to_csc_hs_me1a_even[ 84]     =   8'd170;
	gem_pad_to_csc_hs_me1a_even[ 85]     =   8'd170;
	gem_pad_to_csc_hs_me1a_even[ 86]     =   8'd171;
	gem_pad_to_csc_hs_me1a_even[ 87]     =   8'd171;
	gem_pad_to_csc_hs_me1a_even[ 88]     =   8'd172;
	gem_pad_to_csc_hs_me1a_even[ 89]     =   8'd172;
	gem_pad_to_csc_hs_me1a_even[ 90]     =   8'd173;
	gem_pad_to_csc_hs_me1a_even[ 91]     =   8'd173;
	gem_pad_to_csc_hs_me1a_even[ 92]     =   8'd174;
	gem_pad_to_csc_hs_me1a_even[ 93]     =   8'd174;
	gem_pad_to_csc_hs_me1a_even[ 94]     =   8'd175;
	gem_pad_to_csc_hs_me1a_even[ 95]     =   8'd175;
	gem_pad_to_csc_hs_me1a_even[ 96]     =   8'd176;
	gem_pad_to_csc_hs_me1a_even[ 97]     =   8'd176;
	gem_pad_to_csc_hs_me1a_even[ 98]     =   8'd177;
	gem_pad_to_csc_hs_me1a_even[ 99]     =   8'd177;
	gem_pad_to_csc_hs_me1a_even[100]     =   8'd178;
	gem_pad_to_csc_hs_me1a_even[101]     =   8'd178;
	gem_pad_to_csc_hs_me1a_even[102]     =   8'd179;
	gem_pad_to_csc_hs_me1a_even[103]     =   8'd179;
	gem_pad_to_csc_hs_me1a_even[104]     =   8'd180;
	gem_pad_to_csc_hs_me1a_even[105]     =   8'd180;
	gem_pad_to_csc_hs_me1a_even[106]     =   8'd180;
	gem_pad_to_csc_hs_me1a_even[107]     =   8'd181;
	gem_pad_to_csc_hs_me1a_even[108]     =   8'd181;
	gem_pad_to_csc_hs_me1a_even[109]     =   8'd182;
	gem_pad_to_csc_hs_me1a_even[110]     =   8'd182;
	gem_pad_to_csc_hs_me1a_even[111]     =   8'd183;
	gem_pad_to_csc_hs_me1a_even[112]     =   8'd183;
	gem_pad_to_csc_hs_me1a_even[113]     =   8'd184;
	gem_pad_to_csc_hs_me1a_even[114]     =   8'd184;
	gem_pad_to_csc_hs_me1a_even[115]     =   8'd185;
	gem_pad_to_csc_hs_me1a_even[116]     =   8'd185;
	gem_pad_to_csc_hs_me1a_even[117]     =   8'd186;
	gem_pad_to_csc_hs_me1a_even[118]     =   8'd186;
	gem_pad_to_csc_hs_me1a_even[119]     =   8'd187;
	gem_pad_to_csc_hs_me1a_even[120]     =   8'd187;
	gem_pad_to_csc_hs_me1a_even[121]     =   8'd188;
	gem_pad_to_csc_hs_me1a_even[122]     =   8'd188;
	gem_pad_to_csc_hs_me1a_even[123]     =   8'd189;
	gem_pad_to_csc_hs_me1a_even[124]     =   8'd189;
	gem_pad_to_csc_hs_me1a_even[125]     =   8'd190;
	gem_pad_to_csc_hs_me1a_even[126]     =   8'd190;
	gem_pad_to_csc_hs_me1a_even[127]     =   8'd191;
	gem_pad_to_csc_hs_me1a_even[128]     =   8'd191;
	gem_pad_to_csc_hs_me1a_even[129]     =   8'd191;
	gem_pad_to_csc_hs_me1a_even[130]     =   8'd192;
	gem_pad_to_csc_hs_me1a_even[131]     =   8'd192;
	gem_pad_to_csc_hs_me1a_even[132]     =   8'd193;
	gem_pad_to_csc_hs_me1a_even[133]     =   8'd193;
	gem_pad_to_csc_hs_me1a_even[134]     =   8'd194;
	gem_pad_to_csc_hs_me1a_even[135]     =   8'd194;
	gem_pad_to_csc_hs_me1a_even[136]     =   8'd195;
	gem_pad_to_csc_hs_me1a_even[137]     =   8'd195;
	gem_pad_to_csc_hs_me1a_even[138]     =   8'd196;
	gem_pad_to_csc_hs_me1a_even[139]     =   8'd196;
	gem_pad_to_csc_hs_me1a_even[140]     =   8'd197;
	gem_pad_to_csc_hs_me1a_even[141]     =   8'd197;
	gem_pad_to_csc_hs_me1a_even[142]     =   8'd198;
	gem_pad_to_csc_hs_me1a_even[143]     =   8'd198;
	gem_pad_to_csc_hs_me1a_even[144]     =   8'd199;
	gem_pad_to_csc_hs_me1a_even[145]     =   8'd199;
	gem_pad_to_csc_hs_me1a_even[146]     =   8'd200;
	gem_pad_to_csc_hs_me1a_even[147]     =   8'd200;
	gem_pad_to_csc_hs_me1a_even[148]     =   8'd201;
	gem_pad_to_csc_hs_me1a_even[149]     =   8'd201;
	gem_pad_to_csc_hs_me1a_even[150]     =   8'd201;
	gem_pad_to_csc_hs_me1a_even[151]     =   8'd202;
	gem_pad_to_csc_hs_me1a_even[152]     =   8'd202;
	gem_pad_to_csc_hs_me1a_even[153]     =   8'd203;
	gem_pad_to_csc_hs_me1a_even[154]     =   8'd203;
	gem_pad_to_csc_hs_me1a_even[155]     =   8'd204;
	gem_pad_to_csc_hs_me1a_even[156]     =   8'd204;
	gem_pad_to_csc_hs_me1a_even[157]     =   8'd205;
	gem_pad_to_csc_hs_me1a_even[158]     =   8'd205;
	gem_pad_to_csc_hs_me1a_even[159]     =   8'd206;
	gem_pad_to_csc_hs_me1a_even[160]     =   8'd206;
	gem_pad_to_csc_hs_me1a_even[161]     =   8'd207;
	gem_pad_to_csc_hs_me1a_even[162]     =   8'd207;
	gem_pad_to_csc_hs_me1a_even[163]     =   8'd208;
	gem_pad_to_csc_hs_me1a_even[164]     =   8'd208;
	gem_pad_to_csc_hs_me1a_even[165]     =   8'd209;
	gem_pad_to_csc_hs_me1a_even[166]     =   8'd209;
	gem_pad_to_csc_hs_me1a_even[167]     =   8'd210;
	gem_pad_to_csc_hs_me1a_even[168]     =   8'd210;
	gem_pad_to_csc_hs_me1a_even[169]     =   8'd210;
	gem_pad_to_csc_hs_me1a_even[170]     =   8'd211;
	gem_pad_to_csc_hs_me1a_even[171]     =   8'd211;
	gem_pad_to_csc_hs_me1a_even[172]     =   8'd212;
	gem_pad_to_csc_hs_me1a_even[173]     =   8'd212;
	gem_pad_to_csc_hs_me1a_even[174]     =   8'd213;
	gem_pad_to_csc_hs_me1a_even[175]     =   8'd213;
	gem_pad_to_csc_hs_me1a_even[176]     =   8'd214;
	gem_pad_to_csc_hs_me1a_even[177]     =   8'd214;
	gem_pad_to_csc_hs_me1a_even[178]     =   8'd215;
	gem_pad_to_csc_hs_me1a_even[179]     =   8'd215;
	gem_pad_to_csc_hs_me1a_even[180]     =   8'd216;
	gem_pad_to_csc_hs_me1a_even[181]     =   8'd216;
	gem_pad_to_csc_hs_me1a_even[182]     =   8'd217;
	gem_pad_to_csc_hs_me1a_even[183]     =   8'd217;
	gem_pad_to_csc_hs_me1a_even[184]     =   8'd218;
	gem_pad_to_csc_hs_me1a_even[185]     =   8'd218;
	gem_pad_to_csc_hs_me1a_even[186]     =   8'd219;
	gem_pad_to_csc_hs_me1a_even[187]     =   8'd219;
	gem_pad_to_csc_hs_me1a_even[188]     =   8'd219;
	gem_pad_to_csc_hs_me1a_even[189]     =   8'd220;
	gem_pad_to_csc_hs_me1a_even[190]     =   8'd220;
	gem_pad_to_csc_hs_me1a_even[191]     =   8'd221;
  end

endmodule
