`timescale 1ns / 1ps
//-----------------------------------------------------------------------------------------------------------------------
//
//	Variable depth, single bit SRL16E-based parallel shifter
//
//	06/25/10 Initial
//	09/16/10 Port to ise 12
//	10/05/10 Check non-blocking operator, add reg init
//-----------------------------------------------------------------------------------------------------------------------
	module srl16e_bit(clock,adr,d,q);

//-------------------------------------------------------------------------------------------------------------------
// Generics caller may override
//-------------------------------------------------------------------------------------------------------------------
	parameter ADR_WIDTH = 8;		// Addess width
	parameter SRL_DEPTH = 256;		// Shift register stages may be less than 2**ADR_WIDTH

	initial	$display("srl16e_bit: ADR_WIDTH=%d",ADR_WIDTH);
	initial	$display("srl16e_bit: SRL_DEPTH=%d",SRL_DEPTH);

//-------------------------------------------------------------------------------------------------------------------
// Ports
//-------------------------------------------------------------------------------------------------------------------
	input					clock;
	input	[ADR_WIDTH-1:0]	adr;
	input					d;
	output					q;

// Shift d left by adr places
	reg [SRL_DEPTH-1:0] srl=0;

	always @(posedge clock) begin
	srl <= {srl[SRL_DEPTH-2:0], d};
	end

	assign q = srl[adr];
	
//-----------------------------------------------------------------------------------------------------------------------
	endmodule
//-----------------------------------------------------------------------------------------------------------------------
